library verilog;
use verilog.vl_types.all;
entity FINAL2_vlg_vec_tst is
end FINAL2_vlg_vec_tst;
