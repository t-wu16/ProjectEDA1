library verilog;
use verilog.vl_types.all;
entity FINAL_vlg_vec_tst is
end FINAL_vlg_vec_tst;
